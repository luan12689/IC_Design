module test ()